module mux32to1(d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,
	d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,
	d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,S,Y);
	input wire [7:0]	d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31;
	input wire [5:0]  S;
	output reg [7:0] Y;
	
		always@(*) begin
			case(S)
			5'b00000: Y= d0;
			5'b00001: Y= d1;
			5'b00010: Y= d2;
			5'b00011: Y= d3;
			5'b00100: Y= d4;
			5'b00101: Y= d5;
			5'b00110: Y= d6;
			5'b00111: Y= d7;
			5'b01000: Y= d8;
			5'b01001: Y= d9;
			5'b01010: Y= d10;
			5'b01011: Y= d11;
			5'b01100: Y= d12;
			5'b01101: Y= d13;
			5'b01110: Y= d14;
			5'b01111: Y= d15;
			//
			5'b10000: Y= d16;
			5'b10001: Y= d17;
			5'b10010: Y= d18;
			5'b10011: Y= d19;
			5'b10100: Y= d20;
			5'b10101: Y= d21;
			5'b10110: Y= d22;
			5'b10111: Y= d23;
			5'b11000: Y= d24;
			5'b11001: Y= d25;
			5'b11010: Y= d26;
			5'b11011: Y= d27;
			5'b11100: Y= d28;
			5'b11101: Y= d29;
			5'b11110: Y= d30;
			5'b11111: Y= d31;
			endcase
		end
endmodule
