
module demux1to32(d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,
			d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,
			d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,S,W);
	input wire [7:0] W;
	input wire[5:0] S;
	output reg [7:0] d0,d1,d2,d3,d4,d5,d6,d7,d8,d9,d10,d11,d12,d13,d14,d15,d16,d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31;
	
	always@(*) begin
		case(S)
			5'b00000: d0=W;
			5'b00001: d1=W;
			5'b00010: d2=W;
			5'b00011: d3=W;
			5'b00100: d4=W;
			5'b00101: d5=W;
			5'b00110: d6=W;
			5'b00111: d7=W;
			5'b01000: d8=W;
			5'b01001: d9=W;
			5'b01010: d10=W;
			5'b01011: d11=W;
			5'b01100: d12=W;
			5'b01101: d13=W;
			5'b01110: d14=W;
			5'b01111: d15=W;
			//
			5'b10000: d16=W;
			5'b10001: d17=W;
			5'b10010: d18=W;
			5'b10011: d19=W;
			5'b10100: d20=W;
			5'b10101: d21=W;
			5'b10110: d22=W;
			5'b10111: d23=W;
			5'b11000: d24=W;
			5'b11001: d25=W;
			5'b11010: d26=W;
			5'b11011: d27=W;
			5'b11100: d28=W;
			5'b11101: d29=W;
			5'b11110: d30=W;
			5'b11111: d31=W;
		endcase
	end
endmodule